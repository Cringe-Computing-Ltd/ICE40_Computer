module ice_bram(
    // Read port
    input           rclk,
    input   [7:0]   raddr,
    output  [15:0]  rdata,

    // Write port
    input           wclk,
    input           we,
    input   [7:0]   waddr,
    input   [15:0]  wdata,
);

    SB_RAM40_4K SB_RAM40_4K_inst(
        .RDATA(rdata), .RADDR(raddr), .WADDR(waddr), .MASK(16'h0000), .WDATA(wdata), .RCLKE(1), .RCLK(rclk), .RE(1), .WCLKE(1), .WCLK(wclk), .WE(we)
    );
endmodule

module ice_rom(
    // Read port
    input           rclk,
    input   [7:0]   raddr,
    output  [15:0]  rdata,

    // Write port
    input           wclk,
    input           we,
    input   [7:0]   waddr,
    input   [15:0]  wdata,
);

    SB_RAM40_4K SB_RAM40_4K_inst(
        .RDATA(rdata), .RADDR(raddr), .WADDR(waddr), .MASK(16'h0000), .WDATA(wdata), .RCLKE(1), .RCLK(rclk), .RE(1), .WCLKE(1), .WCLK(wclk), .WE(we)
    );

    defparam SB_RAM40_4K_inst.INIT_0 = 256'h000000000000000000000000000000000800000c0F0000002000000c1E0C0000;
    defparam SB_RAM40_4K_inst.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam SB_RAM40_4K_inst.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
endmodule